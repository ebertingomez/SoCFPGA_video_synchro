`default_nettype none
module mire (
    ports
);
    
endmodule