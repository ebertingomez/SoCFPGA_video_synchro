`default_nettype none
module wshb_intercon (
    ports
);
    
endmodule